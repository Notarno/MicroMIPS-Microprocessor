library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ControlUnit is
	port(Op, Fn: in std_logic_vector(5 downto 0);
		  RegWrite, DataRead, DataWrite, ALUSrc, ADDSUB: out std_logic;
		  RegDst, BrType, RegInSrc, PCSrc, LogicFn, FnClass: out std_logic_vector(1 downto 0));
end entity ControlUnit;

architecture func of ControlUnit is
begin
	process(Op, Fn)
	begin
		if (Op = "000000") then
			if (Fn = "100000") then --Add
				RegWrite <= '1';
				RegDst <= "01";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '0';
				ADDSUB <= '0';
				FnClass <= "10";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
			elsif (Fn = "100010") then --Subtract
				RegWrite <= '1';
				RegDst <= "01";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '0';
				ADDSUB <= '1';
				FnClass <= "10";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
			elsif (Fn = "101010") then --Set Less Than
				RegWrite <= '1';
				RegDst <= "01";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '0';
				ADDSUB <= '1';
				FnClass <= "01";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
			elsif (Fn = "100100") then --AND
				RegWrite <= '1';
				RegDst <= "01";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '0';
				LogicFn <= "00";
				FnClass <= "11";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
			elsif (Fn = "100101") then --OR
				RegWrite <= '1';
				RegDst <= "01";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '0';
				LogicFn <= "01";
				FnClass <= "11";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
			elsif (Fn = "100110") then --XOR
				RegWrite <= '1';
				RegDst <= "01";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '0';
				LogicFn <= "10";
				FnClass <= "11";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
			elsif (Fn = "001000") then --Jump Register
				RegWrite <= '0';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				PCSrc <= "01";
			elsif (Fn = "001100") then --System Call
				RegWrite <= '0';
				RegDst <= "00";
				PCSrc <= "11";
			end if;
		elsif (Op = "001111") then --LUI
			RegWrite <= '1';
			RegDst <= "00";
			RegInSrc <= "01";
			ALUSrc <= '1';
			FnClass <= "00";
			DataRead <= '0';
			DataWrite <= '0';
			Brtype <= "00";
			PCSrc <= "00";
		elsif (Op = "001000") then --Add Immediate
				RegWrite <= '1';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '1';
				ADDSUB <= '0';
				FnClass <= "10";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
		elsif (Op = "001010") then --Set less than immediate
				RegWrite <= '1';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '1';
				ADDSUB <= '1';
				FnClass <= "01";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
		elsif (Op = "001100") then --AND immediate
				RegWrite <= '1';
				RegDst <= "01";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '1';
				LogicFn <= "00";
				FnClass <= "11";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
		elsif (Op = "001101") then --OR immediate
				RegWrite <= '1';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '1';
				LogicFn <= "01";
				FnClass <= "11";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
		elsif (Op = "001110") then --XOR immediate
				RegWrite <= '1';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				ALUSrc <= '1';
				LogicFn <= "10";
				FnClass <= "11";
				BrType <= "00";
				RegInSrc <= "01";
				PCSrc <= "00";
		elsif (Op = "100011") then --Load Word
				RegWrite <= '1';
				RegDst <= "00";
				DataRead <= '1';
				DataWrite <= '0';
				ALUSrc <= '1';
				ADDSUB <= '0';
				FnClass <= "10";
				BrType <= "00";
				RegInSrc <= "00";
				PCSrc <= "00";
		elsif (Op = "101011") then --Store Word
				RegWrite <= '1';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '1';
				ALUSrc <= '1';
				ADDSUB <= '0';
				FnClass <= "10";
				BrType <= "00";
				PCSrc <= "00";
		elsif (Op = "000010") then --Jump
				RegWrite <= '0';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				PCSrc <= "01";
		elsif (Op = "000001") then --Branch on less than 0
				RegWrite <= '0';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				BrType <= "11";
				PCSrc <= "00";
		elsif (Op = "000100") then --Branch on equal
				RegWrite <= '0';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				BrType <= "01";
				PCSrc <= "00";
		elsif (Op = "000101") then --Branch on Not equal
				RegWrite <= '0';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				BrType <= "10";
				PCSrc <= "00";
		elsif (Op = "000011") then --Jump and Link
				RegWrite <= '1';
				RegDst <= "00";
				DataRead <= '0';
				DataWrite <= '0';
				BrType <= "00";
				PCSrc <= "01";
		end if;
	end process;
end architecture func;